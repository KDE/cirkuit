%%backend=circuitmacros%%
\documentclass{article}
\usepackage[utf8x]{inputenc}

\usepackage{pstricks,pst-eps,graphicx,ifpdf,pst-grad,amsmath,wasysym}
\usepackage{sansmath}
\usepackage{lmodern}
\pagestyle{empty}
\thispagestyle{empty}

\begin{document}
\newbox\graph
\sffamily
\sansmath
\begin{TeXtoEPS}
%%SOURCE%%
\box
\graph
\end{TeXtoEPS}
\end{document}

