%%backend=circuitmacros%%
\documentclass{article}
\usepackage[utf8x]{inputenc}
\usepackage{tikz,amsmath}

\usetikzlibrary{arrows,snakes,backgrounds,patterns,matrix,shapes,fit,calc,shadows,plotmarks}
\usepackage[graphics,tightpage,active]{preview}
\PreviewEnvironment{tikzpicture}
\PreviewEnvironment{equation}
\PreviewEnvironment{equation*}
\newlength{\imagewidth}
\newlength{\imagescale}
\pagestyle{empty}

\begin{document}
\thispagestyle{empty}
%%SOURCE%%
\end{document}
