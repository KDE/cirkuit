%%backend=pstricks%%
\documentclass{article}
\usepackage[utf8x]{inputenc}

\usepackage[dvipsnames,svgnames]{pstricks}
\usepackage{pst-eps,graphicx,pst-grad,pst-circ,amsmath}
\usepackage{pst-node}
\usepackage{pst-coil}
\usepackage{pst-ob3d}
\usepackage{pstricks-add}
\usepackage{pst-labo}
\usepackage{pst-optic}
\usepackage{pst-osci}
\usepackage{pst-spectra}
\usepackage{pst-eucl}
\usepackage{pst-bar}
\usepackage{filecontents}
\usepackage{pst-func}
\usepackage{pst-blur}

\pagestyle{empty}
\thispagestyle{empty}

% ppl - palatino
% pbk = bookman
% phv = helvetiva
% cmtt - computer modern
% cmr  - computer modern roman - default
% ptm  - times
% cmss - computer modern san serif
% lmtt - latin modern typewriter
% see: http://www.tug.dk/FontCatalogue/
%
% in texlive-fonts-extra kp and other fonts
%  listing installed files gives internsl names.
%  at present time installing this package causes psfont errors in PyX
% jkpl - kp light
% jkp  - kp
% jkptt - teletype
% jkpss  - san serif

\begin{document}
{\fontfamily{jkpss}\selectfont
\newbox
\graph

\begin{TeXtoEPS}
%%SOURCE%%
\box
\graph
\end{TeXtoEPS}
}
\end{document}

