%%backend=pstricks%%
\documentclass{article}

\usepackage{pstricks,pst-eps,graphicx,pst-grad,amsmath}
\pagestyle{empty}
\thispagestyle{empty}

\begin{document}
\newbox\graph
\begin{TeXtoEPS}
%%SOURCE%%
\box
\graph
\end{TeXtoEPS}
\end{document}