%%backend=tikz%%
%\documentclass{article}
\documentclass[tikz, border=10pt, 12pt]{standalone}

\usepackage{amsmath}
\usepackage{tikz}
\usepackage{verbatim}
\usepackage[europeanresistors,americaninductors,siunitx]{circuitikz}
\usetikzlibrary{arrows,decorations,backgrounds,patterns,matrix,shapes,fit,calc,shadows,plotmarks}
\usepackage[graphics,tightpage,active]{preview}
\usepackage{smartdiagram}

\PreviewEnvironment{tikzpicture}
\PreviewEnvironment{equation}
\PreviewEnvironment{equation*}
\pagestyle{empty}

\begin{document}
\thispagestyle{empty}
%%SOURCE%%
\end{document}
